
interface intf();
    // ------------------- port declaration-------------------------------------
    logic [7:0] in;
    logic [2:0] sel;
    logic       out;
    //--------------------------------------------------------------------------

endinterface

